module name_tb;
reg [4:0]a;
wire y;
name uut(.a(a),.y(y));
initial begin
//M
a=5'b11111;
#5;
a = 5'b11000;
#5;
a = 5'b00100;
#5;
a= 5'b11000;
#5;
a=5'b11111;
#5;
//gap
a=5'b00000;
#5;
//E
a=5'b11111;
#5;
a=5'b10101;
#5;
a=5'b10101;
#5;
a=5'b10001;
#5;
a=5'b10001;
#5;
//gap
a=5'b00000;
#5;
//E
a=5'b11111;
#5;
a=5'b10101;
#5;
a=5'b10101;
#5;
a=5'b10001;
#5;
a=5'b10001;
#5;
//gap
a=5'b00000;
#5;
//N
a=5'b11111;
#5;
a=5'b10000;
#5;
a=5'b11111;
#5;
a=5'b00001;
#5;
a=5'b11111;
#5;
//gap
a=5'b00000;
#5;
//A
a=5'b11111;
#5;
a=5'b10100;
#5;
a=5'b10100;
#5;
a=5'b10100;
#5;
a=5'b11111;
#5;
//gap
a=5'b00000;
#5;
//K
a=5'b11111;
#5;
a=5'b00100;
#5;
a=5'b00100;
#5;
a=5'b01010;
#5;
a=5'b10001;
#5;
//gap
a=5'b00000;
#5;
//S
a=5'b11101;
#5;
a=5'b10101;
#5;
a=5'b10101;
#5;
a=5'b10101;
#5;
a=5'b10111;
#5;
//gap
a=5'b00000;
#5;
//H
a=5'b11111;
#5;
a=5'b00100;
#5;
a=5'b00100;
#5;
a=5'b00100;
#5;
a=5'b11111;
#5;
//gap
a=5'b00000;
#5;
//I
a=5'b10001;
#5;
a=5'b10001;
#5;
a=5'b11111;
#5;
a=5'b10001;
#5;
a=5'b10001;
#5;
//gap
a=5'b00000;
#5;
end 
endmodule
